f := ld_r_r(state, f, r(y), r(z));
